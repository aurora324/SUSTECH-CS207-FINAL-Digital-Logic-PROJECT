`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2024/01/01 10:25:12
// Design Name: 
// Module Name: music_lib
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module music_lib(
    input clk,
    input [4:0] in_note,
    input RorW,
    input back_to_start,
    input [2:0] song_select,
    output reg [4:0] note,
    output[8:0] out_state
    );
    reg[8:0] state = 0;
    reg[8:0] next_state;
    
    wire[4:0] song1 [0:511];
    wire[4:0] song2 [0:511];
    wire[4:0] song3 [0:511];
    wire[4:0] song4 [0:511];
    reg[4:0] song5 [0:511];
    reg[4:0] song6 [0:511];
    reg[4:0] song7 [0:511];
    reg[4:0] song8 [0:511];
    
    assign song1[511] = 5'b11111;
    assign song2[511] = 5'b11111;
    assign song3[511] = 5'b11111;
    assign song4[511] = 5'b11111;
    
    assign song1[0]=5'b0_0001;
    assign song1[1]=5'b0_0001;
    assign song1[2]=5'b0_0000;
    assign song1[3]=5'b0_0000;
    assign song1[4]=5'b0_0001;
    assign song1[5]=5'b0_0001;
    assign song1[6]=5'b0_0000;
    assign song1[7]=5'b0_0000;
    assign song1[8]=5'b0_0101;
    assign song1[9]=5'b0_0101;
    assign song1[10]=5'b0_0000;
    assign song1[11]=5'b0_0000;
    assign song1[12]=5'b0_0101;
    assign song1[13]=5'b0_0101;
    assign song1[14]=5'b0_0000;
    assign song1[15]=5'b0_0000;
    assign song1[16]=5'b0_0110;
    assign song1[17]=5'b0_0110;
    assign song1[18]=5'b0_0000;
    assign song1[19]=5'b0_0000;
    assign song1[20]=5'b0_0110;
    assign song1[21]=5'b0_0110;
    assign song1[22]=5'b0_0000;
    assign song1[23]=5'b0_0000;
    assign song1[24]=5'b0_0101;
    assign song1[25]=5'b0_0101;
    assign song1[26]=5'b0_0000;
    assign song1[27]=5'b0_0000;
    assign song1[28]=5'b0_0100;
    assign song1[29]=5'b0_0100;
    assign song1[30]=5'b0_0000;
    assign song1[31]=5'b0_0000;
    assign song1[32]=5'b0_0100;
    assign song1[33]=5'b0_0100;
    assign song1[34]=5'b0_0000;
    assign song1[35]=5'b0_0000;
    assign song1[36]=5'b0_0011;
    assign song1[37]=5'b0_0011;
    assign song1[38]=5'b0_0000;
    assign song1[39]=5'b0_0000;
    assign song1[40]=5'b0_0011;
    assign song1[41]=5'b0_0011;
    assign song1[42]=5'b0_0000;
    assign song1[43]=5'b0_0000;
    assign song1[44]=5'b0_0010;
    assign song1[45]=5'b0_0010;
    assign song1[46]=5'b0_0000;
    assign song1[47]=5'b0_0000;
    assign song1[48]=5'b0_0010;
    assign song1[49]=5'b0_0010;
    assign song1[50]=5'b0_0000;
    assign song1[51]=5'b0_0000;
    assign song1[52]=5'b0_0001;
    assign song1[53]=5'b0_0001;
    assign song1[54]=5'b0_0000;
    assign song1[55]=5'b0_0000;
    assign song1[56]=5'b0_0101;
    assign song1[57]=5'b0_0101;
    assign song1[58]=5'b0_0000;
    assign song1[59]=5'b0_0000;
    assign song1[60]=5'b0_0101;
    assign song1[61]=5'b0_0101;
    assign song1[62]=5'b0_0000;
    assign song1[63]=5'b0_0000;
    assign song1[64]=5'b0_0100;
    assign song1[65]=5'b0_0100;
    assign song1[66]=5'b0_0000;
    assign song1[67]=5'b0_0000;
    assign song1[68]=5'b0_0100;
    assign song1[69]=5'b0_0100;
    assign song1[70]=5'b0_0000;
    assign song1[71]=5'b0_0000;
    assign song1[72]=5'b0_0011;
    assign song1[73]=5'b0_0011;
    assign song1[74]=5'b0_0000;
    assign song1[75]=5'b0_0000;
    assign song1[76]=5'b0_0011;
    assign song1[77]=5'b0_0011;
    assign song1[78]=5'b0_0000;
    assign song1[79]=5'b0_0000;
    assign song1[80]=5'b0_0010;
    assign song1[81]=5'b0_0010;
    assign song1[82]=5'b0_0000;
    assign song1[83]=5'b0_0000;
    assign song1[84]=5'b0_0101;
    assign song1[85]=5'b0_0101;
    assign song1[86]=5'b0_0000;
    assign song1[87]=5'b0_0000;
    assign song1[88]=5'b0_0101;
    assign song1[89]=5'b0_0101;
    assign song1[90]=5'b0_0000;
    assign song1[91]=5'b0_0000;
    assign song1[92]=5'b0_0100;
    assign song1[93]=5'b0_0100;
    assign song1[94]=5'b0_0000;
    assign song1[95]=5'b0_0000;
    assign song1[96]=5'b0_0100;
    assign song1[97]=5'b0_0100;
    assign song1[98]=5'b0_0000;
    assign song1[99]=5'b0_0000;
    assign song1[100]=5'b0_0011;
    assign song1[101]=5'b0_0011;
    assign song1[102]=5'b0_0000;
    assign song1[103]=5'b0_0000;
    assign song1[104]=5'b0_0011;
    assign song1[105]=5'b0_0011;
    assign song1[106]=5'b0_0000;
    assign song1[107]=5'b0_0000;
    assign song1[108]=5'b0_0010;
    assign song1[109]=5'b0_0010;
    assign song1[110]=5'b0_0000;
    assign song1[111]=5'b0_0000;
    assign song1[112]=5'b0_0001;
    assign song1[113]=5'b0_0001;
    assign song1[114]=5'b0_0000;
    assign song1[115]=5'b0_0000;
    assign song1[116]=5'b0_0001;
    assign song1[117]=5'b0_0001;
    assign song1[118]=5'b0_0000;
    assign song1[119]=5'b0_0000;
    assign song1[120]=5'b0_0101;
    assign song1[121]=5'b0_0101;
    assign song1[122]=5'b0_0000;
    assign song1[123]=5'b0_0000;
    assign song1[124]=5'b0_0101;
    assign song1[125]=5'b0_0101;
    assign song1[126]=5'b0_0000;
    assign song1[127]=5'b0_0000;
    assign song1[128]=5'b0_0110;
    assign song1[129]=5'b0_0110;
    assign song1[130]=5'b0_0000;
    assign song1[131]=5'b0_0000;
    assign song1[132]=5'b0_0110;
    assign song1[133]=5'b0_0110;
    assign song1[134]=5'b0_0000;
    assign song1[135]=5'b0_0000;
    assign song1[136]=5'b0_0101;
    assign song1[137]=5'b0_0101;
    assign song1[138]=5'b0_0000;
    assign song1[139]=5'b0_0000;
    assign song1[140]=5'b0_0100;
    assign song1[141]=5'b0_0100;
    assign song1[142]=5'b0_0000;
    assign song1[143]=5'b0_0000;
    assign song1[144]=5'b0_0100;
    assign song1[145]=5'b0_0100;
    assign song1[146]=5'b0_0000;
    assign song1[147]=5'b0_0000;
    assign song1[148]=5'b0_0011;
    assign song1[149]=5'b0_0011;
    assign song1[150]=5'b0_0000;
    assign song1[151]=5'b0_0000;
    assign song1[152]=5'b0_0011;
    assign song1[153]=5'b0_0011;
    assign song1[154]=5'b0_0000;
    assign song1[155]=5'b0_0000;
    assign song1[156]=5'b0_0010;
    assign song1[157]=5'b0_0010;
    assign song1[158]=5'b0_0000;
    assign song1[159]=5'b0_0000;
    assign song1[160]=5'b0_0010;
    assign song1[161]=5'b0_0010;
    assign song1[162]=5'b0_0000;
    assign song1[163]=5'b0_0000;
    assign song1[164]=5'b0_0001;
    assign song1[165]=5'b0_0001;
    assign song1[166]=5'b0_0000;
    assign song1[167]=5'b0_0000;
    assign song1[168]=5'd31  ;

assign  song2[0]=5'd5  ;
assign  song2[1]=5'd0  ;
assign  song2[2]=5'd5  ;
assign  song2[3]=5'd0  ;
assign  song2[4]=5'd15  ;
assign  song2[5]=5'd15  ;
assign  song2[6]=5'd0  ;
assign  song2[7]=5'd0  ;
assign  song2[8]=5'd15  ;
assign  song2[9]=5'd0  ;
assign  song2[10]=5'd16  ;
assign  song2[11]=5'd0  ;
assign  song2[12]=5'd15  ;
assign  song2[13]=5'd0  ;
assign  song2[14]=5'd7  ;
assign  song2[15]=5'd0  ;
assign  song2[16]=5'd6  ;
assign  song2[17]=5'd6  ;
assign  song2[18]=5'd0  ;
assign  song2[19]=5'd0  ;
assign  song2[20]=5'd6  ;
assign  song2[21]=5'd6  ;
assign  song2[22]=5'd0  ;
assign  song2[23]=5'd0  ;
assign  song2[24]=5'd6  ;
assign  song2[25]=5'd0  ;
assign  song2[26]=5'd6  ;
assign  song2[27]=5'd0  ;
assign  song2[28]=5'd16  ;
assign  song2[29]=5'd16  ;
assign  song2[30]=5'd0  ;
assign  song2[31]=5'd0  ;
assign  song2[32]=5'd16  ;
assign  song2[33]=5'd0  ;
assign  song2[34]=5'd17  ;
assign  song2[35]=5'd0  ;
assign  song2[36]=5'd16  ;
assign  song2[37]=5'd0  ;
assign  song2[38]=5'd15  ;
assign  song2[39]=5'd0  ;
assign  song2[40]=5'd7  ;
assign  song2[41]=5'd7  ;
assign  song2[42]=5'd0  ;
assign  song2[43]=5'd0  ;
assign  song2[44]=5'd5  ;
assign  song2[45]=5'd5  ;
assign  song2[46]=5'd0  ;
assign  song2[47]=5'd0  ;
assign  song2[48]=5'd5  ;
assign  song2[49]=5'd0  ;
assign  song2[50]=5'd5  ;
assign  song2[51]=5'd0  ;
assign  song2[52]=5'd17  ;
assign  song2[53]=5'd17  ;
assign  song2[54]=5'd0  ;
assign  song2[55]=5'd0  ;
assign  song2[56]=5'd17  ;
assign  song2[57]=5'd0  ;
assign  song2[58]=5'd18  ;
assign  song2[59]=5'd0  ;
assign  song2[60]=5'd17  ;
assign  song2[61]=5'd0  ;
assign  song2[62]=5'd16  ;
assign  song2[63]=5'd0  ;
assign  song2[64]=5'd15  ;
assign  song2[65]=5'd15  ;
assign  song2[66]=5'd0  ;
assign  song2[67]=5'd0  ;
assign  song2[68]=5'd6  ;
assign  song2[69]=5'd6  ;
assign  song2[70]=5'd0  ;
assign  song2[71]=5'd0  ;
assign  song2[72]=5'd5  ;
assign  song2[73]=5'd0  ;
assign  song2[74]=5'd5  ;
assign  song2[75]=5'd0  ;
assign  song2[76]=5'd6  ;
assign  song2[77]=5'd6  ;
assign  song2[78]=5'd0  ;
assign  song2[79]=5'd0  ;
assign  song2[80]=5'd16  ;
assign  song2[81]=5'd16  ;
assign  song2[82]=5'd0  ;
assign  song2[83]=5'd0  ;
assign  song2[84]=5'd7  ;
assign  song2[85]=5'd7  ;
assign  song2[86]=5'd0  ;
assign  song2[87]=5'd0  ;
assign  song2[88]=5'd15  ;
assign  song2[89]=5'd15  ;
assign  song2[90]=5'd15  ;
assign  song2[91]=5'd15  ;
assign  song2[92]=5'd0  ;
assign  song2[93]=5'd0  ;
assign  song2[94]=5'd5  ;
assign  song2[95]=5'd0  ;
assign  song2[96]=5'd5  ;
assign  song2[97]=5'd0  ;
assign  song2[98]=5'd15  ;
assign  song2[99]=5'd15  ;
assign  song2[100]=5'd0  ;
assign  song2[101]=5'd0  ;
assign  song2[102]=5'd15  ;
assign  song2[103]=5'd15  ;
assign  song2[104]=5'd0  ;
assign  song2[105]=5'd0  ;
assign  song2[106]=5'd15  ;
assign  song2[107]=5'd15  ;
assign  song2[108]=5'd0  ;
assign  song2[109]=5'd0  ;
assign  song2[110]=5'd7  ;
assign  song2[111]=5'd7  ;
assign  song2[112]=5'd7  ;
assign  song2[113]=5'd7  ;
assign  song2[114]=5'd0  ;
assign  song2[115]=5'd0  ;
assign  song2[116]=5'd7  ;
assign  song2[117]=5'd0  ;
assign  song2[118]=5'd7  ;
assign  song2[119]=5'd0  ;
assign  song2[120]=5'd15  ;
assign  song2[121]=5'd15  ;
assign  song2[122]=5'd0  ;
assign  song2[123]=5'd0  ;
assign  song2[124]=5'd7  ;
assign  song2[125]=5'd7  ;
assign  song2[126]=5'd0  ;
assign  song2[127]=5'd0  ;
assign  song2[128]=5'd6  ;
assign  song2[129]=5'd6  ;
assign  song2[130]=5'd0  ;
assign  song2[131]=5'd0  ;
assign  song2[132]=5'd5  ;
assign  song2[133]=5'd5  ;
assign  song2[134]=5'd5  ;
assign  song2[135]=5'd5  ;
assign  song2[136]=5'd0  ;
assign  song2[137]=5'd0  ;
assign  song2[138]=5'd16  ;
assign  song2[139]=5'd0  ;
assign  song2[140]=5'd16  ;
assign  song2[141]=5'd0  ;
assign  song2[142]=5'd17  ;
assign  song2[143]=5'd17  ;
assign  song2[144]=5'd0  ;
assign  song2[145]=5'd0  ;
assign  song2[146]=5'd16  ;
assign  song2[147]=5'd16  ;
assign  song2[148]=5'd0  ;
assign  song2[149]=5'd0  ;
assign  song2[150]=5'd15  ;
assign  song2[151]=5'd15  ;
assign  song2[152]=5'd0  ;
assign  song2[153]=5'd0  ;
assign  song2[154]=5'd19  ;
assign  song2[155]=5'd19  ;
assign  song2[156]=5'd0  ;
assign  song2[157]=5'd0  ;
assign  song2[158]=5'd5  ;
assign  song2[159]=5'd5  ;
assign  song2[160]=5'd0  ;
assign  song2[161]=5'd0  ;
assign  song2[162]=5'd5  ;
assign  song2[163]=5'd0  ;
assign  song2[164]=5'd5  ;
assign  song2[165]=5'd0  ;
assign  song2[166]=5'd6  ;
assign  song2[167]=5'd6  ;
assign  song2[168]=5'd0  ;
assign  song2[169]=5'd0  ;
assign  song2[170]=5'd16  ;
assign  song2[171]=5'd16  ;
assign  song2[172]=5'd0  ;
assign  song2[173]=5'd0  ;
assign  song2[174]=5'd7  ;
assign  song2[175]=5'd7  ;
assign  song2[176]=5'd0  ;
assign  song2[177]=5'd0  ;
assign  song2[178]=5'd15  ;
assign  song2[179]=5'd15  ;
assign  song2[180]=5'd15  ;
assign  song2[181]=5'd15  ;
assign  song2[182]=5'd15  ;
assign  song2[183]=5'd15  ;
assign  song2[184]=5'd15  ;
assign  song2[185]=5'd15  ;
assign  song2[186]=5'd31  ;

assign song3[0]=5'd12 ;
assign song3[1]=5'd0 ;
assign song3[2]=5'd12 ;
assign song3[3]=5'd0 ;
assign song3[4]=5'd13 ;
assign song3[5]=5'd13 ;
assign song3[6]=5'd0 ;
assign song3[7]=5'd0 ;
assign song3[8]=5'd12 ;
assign song3[9]=5'd12 ;
assign song3[10]=5'd0 ;
assign song3[11]=5'd0 ;
assign song3[12]=5'd1 ;
assign song3[13]=5'd1 ;
assign song3[14]=5'd0 ;
assign song3[15]=5'd0 ;
assign song3[16]=5'd14 ;
assign song3[17]=5'd14 ;
assign song3[18]=5'd0 ;
assign song3[19]=5'd0 ;
assign song3[20]=5'd12 ;
assign song3[21]=5'd0 ;
assign song3[22]=5'd12 ;
assign song3[23]=5'd0 ;
assign song3[24]=5'd13 ;
assign song3[25]=5'd13 ;
assign song3[26]=5'd0 ;
assign song3[27]=5'd0 ;
assign song3[28]=5'd12 ;
assign song3[29]=5'd12 ;
assign song3[30]=5'd0 ;
assign song3[31]=5'd0 ;
assign song3[32]=5'd2 ;
assign song3[33]=5'd2 ;
assign song3[34]=5'd0 ;
assign song3[35]=5'd0 ;
assign song3[36]=5'd1 ;
assign song3[37]=5'd1 ;
assign song3[38]=5'd0 ;
assign song3[39]=5'd0 ;
assign song3[40]=5'd12 ;
assign song3[41]=5'd12 ;
assign song3[42]=5'd0 ;
assign song3[43]=5'd0 ;
assign song3[44]=5'd12 ;
assign song3[45]=5'd12 ;
assign song3[46]=5'd0 ;
assign song3[47]=5'd0 ;
assign song3[48]=5'd5 ;
assign song3[49]=5'd5 ;
assign song3[50]=5'd0 ;
assign song3[51]=5'd0 ;
assign song3[52]=5'd3 ;
assign song3[53]=5'd3 ;
assign song3[54]=5'd0 ;
assign song3[55]=5'd0 ;
assign song3[56]=5'd1 ;
assign song3[57]=5'd1 ;
assign song3[58]=5'd0 ;
assign song3[59]=5'd0 ;
assign song3[60]=5'd14 ;
assign song3[61]=5'd14 ;
assign song3[62]=5'd0 ;
assign song3[63]=5'd0 ;
assign song3[64]=5'd6 ;
assign song3[65]=5'd6 ;
assign song3[66]=5'd0 ;
assign song3[67]=5'd0 ;
assign song3[68]=5'd4 ;
assign song3[69]=5'd4 ;
assign song3[70]=5'd4 ;
assign song3[71]=5'd0 ;
assign song3[72]=5'd4 ;
assign song3[73]=5'd0 ;
assign song3[74]=5'd3 ;
assign song3[75]=5'd3 ;
assign song3[76]=5'd0 ;
assign song3[77]=5'd0 ;
assign song3[78]=5'd1 ;
assign song3[79]=5'd1 ;
assign song3[80]=5'd0 ;
assign song3[81]=5'd0 ;
assign song3[82]=5'd2 ;
assign song3[83]=5'd2 ;
assign song3[84]=5'd0 ;
assign song3[85]=5'd0 ;
assign song3[86]=5'd1 ;
assign song3[87]=5'd1 ;
assign song3[88]=5'd31 ;

assign song4[0]=5'd20 ;
assign song4[1]=5'd20 ;
assign song4[2]=5'd0 ;
assign song4[3]=5'd0 ;
assign song4[4]=5'd20 ;
assign song4[5]=5'd0 ;
assign song4[6]=5'd20 ;
assign song4[7]=5'd0 ;
assign song4[8]=5'd19 ;
assign song4[9]=5'd19 ;
assign song4[10]=5'd0 ;
assign song4[11]=5'd0 ;
assign song4[12]=5'd19 ;
assign song4[13]=5'd19 ;
assign song4[14]=5'd0 ;
assign song4[15]=5'd0 ;
assign song4[16]=5'd17 ;
assign song4[17]=5'd17 ;
assign song4[18]=5'd0 ;
assign song4[19]=5'd0 ;
assign song4[20]=5'd17 ;
assign song4[21]=5'd17 ;
assign song4[22]=5'd0 ;
assign song4[23]=5'd0 ;
assign song4[24]=5'd15 ;
assign song4[25]=5'd15 ;
assign song4[26]=5'd15 ;
assign song4[27]=5'd15 ;
assign song4[28]=5'd15 ;
assign song4[29]=5'd15 ;
assign song4[30]=5'd0 ;
assign song4[31]=5'd0 ;
assign song4[32]=5'd16 ;
assign song4[33]=5'd0 ;
assign song4[34]=5'd17 ;
assign song4[35]=5'd0 ;
assign song4[36]=5'd16 ;
assign song4[37]=5'd0 ;
assign song4[38]=5'd15 ;
assign song4[39]=5'd0 ;
assign song4[40]=5'd6 ;
assign song4[41]=5'd6 ;
assign song4[42]=5'd0 ;
assign song4[43]=5'd0 ;
assign song4[44]=5'd15 ;
assign song4[45]=5'd15 ;
assign song4[46]=5'd0 ;
assign song4[47]=5'd0 ;
assign song4[48]=5'd6 ;
assign song4[49]=5'd6 ;
assign song4[50]=5'd6 ;
assign song4[51]=5'd6 ;
assign song4[52]=5'd6 ;
assign song4[53]=5'd6 ;
assign song4[54]=5'd0 ;
assign song4[55]=5'd0 ;
assign song4[56]=5'd0 ;
assign song4[57]=5'd0 ;
assign song4[58]=5'd0 ;
assign song4[59]=5'd0 ;
assign song4[60]=5'd0 ;
assign song4[61]=5'd0 ;
assign song4[62]=5'd0 ;
assign song4[63]=5'd0 ;
assign song4[64]=5'd13 ;
assign song4[65]=5'd13 ;
assign song4[66]=5'd0 ;
assign song4[67]=5'd0 ;
assign song4[68]=5'd13 ;
assign song4[69]=5'd0 ;
assign song4[70]=5'd13 ;
assign song4[71]=5'd0 ;
assign song4[72]=5'd2 ;
assign song4[73]=5'd2 ;
assign song4[74]=5'd0 ;
assign song4[75]=5'd0 ;
assign song4[76]=5'd3 ;
assign song4[77]=5'd3 ;
assign song4[78]=5'd0 ;
assign song4[79]=5'd0 ;
assign song4[80]=5'd13 ;
assign song4[81]=5'd13 ;
assign song4[82]=5'd0 ;
assign song4[83]=5'd0 ;
assign song4[84]=5'd13 ;
assign song4[85]=5'd0 ;
assign song4[86]=5'd13 ;
assign song4[87]=5'd0 ;
assign song4[88]=5'd2 ;
assign song4[89]=5'd2 ;
assign song4[90]=5'd0 ;
assign song4[91]=5'd0 ;
assign song4[92]=5'd3 ;
assign song4[93]=5'd3 ;
assign song4[94]=5'd0 ;
assign song4[95]=5'd0 ;
assign song4[96]=5'd17 ;
assign song4[97]=5'd17 ;
assign song4[98]=5'd0 ;
assign song4[99]=5'd0 ;
assign song4[100]=5'd17 ;
assign song4[101]=5'd0 ;
assign song4[102]=5'd16 ;
assign song4[103]=5'd0 ;
assign song4[104]=5'd17 ;
assign song4[105]=5'd17 ;
assign song4[106]=5'd0 ;
assign song4[107]=5'd0 ;
assign song4[108]=5'd19 ;
assign song4[109]=5'd19 ;
assign song4[110]=5'd0 ;
assign song4[111]=5'd0 ;
assign song4[112]=5'd17 ;
assign song4[113]=5'd17 ;
assign song4[114]=5'd17 ;
assign song4[115]=5'd17 ;
assign song4[116]=5'd17 ;
assign song4[117]=5'd17 ;
assign song4[118]=5'd0 ;
assign song4[119]=5'd0 ;
assign song4[120]=5'd15 ;
assign song4[121]=5'd15 ;
assign song4[122]=5'd15 ;
assign song4[123]=5'd15 ;
assign song4[124]=5'd15 ;
assign song4[125]=5'd15 ;
assign song4[126]=5'd0 ;
assign song4[127]=5'd0 ;
assign song4[128]=5'd16 ;
assign song4[129]=5'd0 ;
assign song4[130]=5'd17 ;
assign song4[131]=5'd0 ;
assign song4[132]=5'd16 ;
assign song4[133]=5'd0 ;
assign song4[134]=5'd15 ;
assign song4[135]=5'd0 ;
assign song4[136]=5'd6 ;
assign song4[137]=5'd6 ;
assign song4[138]=5'd0 ;
assign song4[139]=5'd0 ;
assign song4[140]=5'd15 ;
assign song4[141]=5'd15 ;
assign song4[142]=5'd0 ;
assign song4[143]=5'd0 ;
assign song4[144]=5'd17 ;
assign song4[145]=5'd17 ;
assign song4[146]=5'd17 ;
assign song4[147]=5'd0 ;
assign song4[148]=5'd0 ;
assign song4[149]=5'd0 ;
assign song4[150]=5'd16 ;
assign song4[151]=5'd0 ;
assign song4[152]=5'd17 ;
assign song4[153]=5'd17 ;
assign song4[154]=5'd17 ;
assign song4[155]=5'd17 ;
assign song4[156]=5'd17 ;
assign song4[157]=5'd17 ;
assign song4[158]=5'd0 ;
assign song4[159]=5'd0 ;
assign song4[160]=5'd31 ;

    always@(posedge clk,negedge back_to_start)
    begin
    if(!back_to_start)
    begin
        state <= 0;
    end
    else
        state <= next_state;
    end
    //RorW=0 read, RorW=1 write
    always@*
    begin
    next_state = state+1;
    if(RorW)
        begin
        case(song_select)
        3'b100:song5[state] = in_note;
        3'b101:song6[state] = in_note;
        3'b110:song7[state] = in_note;
        3'b111:song8[state] = in_note;
        endcase
        end
    end
    
    always@*
    begin
    if(!back_to_start)
    note = 5'b0_0000;
    else
    begin
    case(song_select)
    3'b000:note = song1[state];
    3'b001:note = song2[state];
    3'b010:note = song3[state];
    3'b011:note = song4[state];
    3'b100:note = song5[state];
    3'b101:note = song6[state];
    3'b110:note = song7[state];
    3'b111:note = song8[state];
    endcase
    end
    end
    
    assign  out_state = state;
endmodule
